/* file: top.v
 Description: Top module for the whole project design with CPU, GPU, NPU, memory, and ILA components
 Author: Jeremy Cai
 Date: Feb. 13, 2026
 Version: 1.0
 */