/* file: fu.v
 Description: Forwarding unit module for the pipeline CPU design
 Author: Jeremy Cai
 Date: Feb. 16, 2026
 Version: 1.0
 */

`ifndef FU_V
`define FU_V

`include "define.v"

`endif // FU_V
