/* file: hdu.v
 Description: Hazard detection unit module for the Arm pipeline CPU design
 Author: Jeremy Cai
 Date: Feb. 16, 2026
 Version: 1.0
 */

`ifndef HDU_V
`define HDU_V

`include "define.v"

`endif // HDU_V
