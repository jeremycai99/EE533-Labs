`ifndef TOP_V
`define TOP_V

`include "define.v"

`include "i_mem.v"
`include "d_mem.v"
`include "cpu.v"

module top (
    input wire clk,
    input wire rst_n
);

// Instantiate instruction memory



`endif // TOP_V
